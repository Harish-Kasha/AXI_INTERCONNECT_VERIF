`define CORE0_OFFSET                     'h000
`define CORE1_OFFSET                     'h800

`define CH0_OFFSET                       'h000
`define CH1_OFFSET                       'h100
`define CH2_OFFSET                       'h200
`define CH3_OFFSET                       'h300
`define CH4_OFFSET                       'h400
`define CH5_OFFSET                       'h500
`define CH6_OFFSET                       'h600
`define CH7_OFFSET                       'h700


`define CMD_REG0_OFFSET                  'h00
`define CMD_REG1_OFFSET                  'h04
`define CMD_REG2_OFFSET                  'h08
`define CMD_REG3_OFFSET                  'h0C
`define STATIC_REG0_OFFSET               'h10
`define STATIC_REG1_OFFSET               'h14
`define STATIC_REG2_OFFSET               'h18
`define STATIC_REG3_OFFSET               'h1C
`define STATIC_REG4_OFFSET               'h20

`define RESTRICT_REG_OFFSET              'h2C
`define READ_OFFSET_REG_OFFSET           'h30
`define WRITE_OFFSET_REG_OFFSET          'h34
`define FIFO_FULLNESS_REG_OFFSET         'h38
`define CMD_OUTS_REG_OFFSET              'h3C
`define CH_ENABLE_REG_OFFSET             'h40
`define CH_START_REG_OFFSET              'h44
`define CH_ACTIVE_REG_OFFSET             'h48
`define COUNT_REG_OFFSET                 'h50
`define INT_RAWSTAT_REG_OFFSET           'hA0
`define INT_CLEAR_REG_OFFSET             'hA4
`define INT_ENABLE_REG_OFFSET            'hA8

`define INT_STATUS_REG_OFFSET            'hAC

`define INT0_STATUS_OFFSET               'h1000

`define CORE0_JOINT_MODE_OFFSET          'h1030
`define CORE1_JOINT_MODE_OFFSET          'h1034

`define CORE0_PRIORITY_OFFSET            'h1038
`define CORE1_PRIORITY_OFFSET            'h103C

`define CORE0_CLKDIV_OFFSET              'h1040
`define CORE1_CLKDIV_OFFSET              'h1044

`define CORE0_CH_START_OFFSET            'h1048
`define CORE1_CH_START_OFFSET            'h104C

`define PERIPH_RX_CTRL_OFFSET            'h1050
`define PERIPH_TX_CTRL_OFFSET            'h1054

`define IDLE_OFFSET                      'h10D0

`define USER_DEF_STATUS_OFFSET           'h10E0

`define USER_CORE0_DEF_STATUS0           'h10F0
`define USER_CORE1_DEF_STATUS0           'h10F8

`define USER_CORE0_DEF_STATUS1           'h10F4
`define USER_CORE1_DEF_STATUS1           'h10FC


