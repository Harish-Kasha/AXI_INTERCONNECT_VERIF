package DMA_rtl_pkg;
  localparam int CMD_REG0_BYTE_WIDTH = 4;
  localparam int CMD_REG0_BYTE_SIZE = 4;
  localparam bit [12:0] CMD_REG0_BYTE_OFFSET = 13'h0000;
  localparam int CMD_REG0_RD_START_ADDR_BIT_WIDTH = 32;
  localparam bit [31:0] CMD_REG0_RD_START_ADDR_BIT_MASK = 32'hffffffff;
  localparam int CMD_REG0_RD_START_ADDR_BIT_OFFSET = 0;
  localparam int CMD_REG1_BYTE_WIDTH = 4;
  localparam int CMD_REG1_BYTE_SIZE = 4;
  localparam bit [12:0] CMD_REG1_BYTE_OFFSET = 13'h0004;
  localparam int CMD_REG1_WR_START_ADDR_BIT_WIDTH = 32;
  localparam bit [31:0] CMD_REG1_WR_START_ADDR_BIT_MASK = 32'hffffffff;
  localparam int CMD_REG1_WR_START_ADDR_BIT_OFFSET = 0;
  localparam int CMD_REG2_BYTE_WIDTH = 4;
  localparam int CMD_REG2_BYTE_SIZE = 4;
  localparam bit [12:0] CMD_REG2_BYTE_OFFSET = 13'h0008;
  localparam int CMD_REG2_BUFFER_SIZE_BIT_WIDTH = 16;
  localparam bit [15:0] CMD_REG2_BUFFER_SIZE_BIT_MASK = 16'hffff;
  localparam int CMD_REG2_BUFFER_SIZE_BIT_OFFSET = 0;
  localparam int CMD_REG3_BYTE_WIDTH = 4;
  localparam int CMD_REG3_BYTE_SIZE = 4;
  localparam bit [12:0] CMD_REG3_BYTE_OFFSET = 13'h000c;
  localparam int CMD_REG3_CMD_SET_INT_BIT_WIDTH = 1;
  localparam bit CMD_REG3_CMD_SET_INT_BIT_MASK = 1'h1;
  localparam int CMD_REG3_CMD_SET_INT_BIT_OFFSET = 0;
  localparam int CMD_REG3_CMD_LAST_BIT_WIDTH = 1;
  localparam bit CMD_REG3_CMD_LAST_BIT_MASK = 1'h1;
  localparam int CMD_REG3_CMD_LAST_BIT_OFFSET = 1;
  localparam int CMD_REG3_CMD_NEXT_ADDR_BIT_WIDTH = 28;
  localparam bit [27:0] CMD_REG3_CMD_NEXT_ADDR_BIT_MASK = 28'hfffffff;
  localparam int CMD_REG3_CMD_NEXT_ADDR_BIT_OFFSET = 4;
  localparam int STATIC_REG0_BYTE_WIDTH = 4;
  localparam int STATIC_REG0_BYTE_SIZE = 4;
  localparam bit [12:0] STATIC_REG0_BYTE_OFFSET = 13'h0010;
  localparam int STATIC_REG0_RD_BURST_MAX_SIZE_BIT_WIDTH = 10;
  localparam bit [9:0] STATIC_REG0_RD_BURST_MAX_SIZE_BIT_MASK = 10'h3ff;
  localparam int STATIC_REG0_RD_BURST_MAX_SIZE_BIT_OFFSET = 0;
  localparam int STATIC_REG0_RD_ALLOW_FULL_BURST_BIT_WIDTH = 1;
  localparam bit STATIC_REG0_RD_ALLOW_FULL_BURST_BIT_MASK = 1'h1;
  localparam int STATIC_REG0_RD_ALLOW_FULL_BURST_BIT_OFFSET = 12;
  localparam int STATIC_REG0_RD_ALLOW_FULL_FIFO_BIT_WIDTH = 1;
  localparam bit STATIC_REG0_RD_ALLOW_FULL_FIFO_BIT_MASK = 1'h1;
  localparam int STATIC_REG0_RD_ALLOW_FULL_FIFO_BIT_OFFSET = 13;
  localparam int STATIC_REG0_RD_TOKENS_BIT_WIDTH = 6;
  localparam bit [5:0] STATIC_REG0_RD_TOKENS_BIT_MASK = 6'h3f;
  localparam int STATIC_REG0_RD_TOKENS_BIT_OFFSET = 16;
  localparam int STATIC_REG0_RD_OUTS_MAX_BIT_WIDTH = 4;
  localparam bit [3:0] STATIC_REG0_RD_OUTS_MAX_BIT_MASK = 4'hf;
  localparam int STATIC_REG0_RD_OUTS_MAX_BIT_OFFSET = 24;
  localparam int STATIC_REG0_RD_OUTSTANDING_BIT_WIDTH = 1;
  localparam bit STATIC_REG0_RD_OUTSTANDING_BIT_MASK = 1'h1;
  localparam int STATIC_REG0_RD_OUTSTANDING_BIT_OFFSET = 30;
  localparam int STATIC_REG0_RD_INCR_BIT_WIDTH = 1;
  localparam bit STATIC_REG0_RD_INCR_BIT_MASK = 1'h1;
  localparam int STATIC_REG0_RD_INCR_BIT_OFFSET = 31;
  localparam int STATIC_REG1_BYTE_WIDTH = 4;
  localparam int STATIC_REG1_BYTE_SIZE = 4;
  localparam bit [12:0] STATIC_REG1_BYTE_OFFSET = 13'h0014;
  localparam int STATIC_REG1_RD_BURST_MAX_SIZE_BIT_WIDTH = 10;
  localparam bit [9:0] STATIC_REG1_RD_BURST_MAX_SIZE_BIT_MASK = 10'h3ff;
  localparam int STATIC_REG1_RD_BURST_MAX_SIZE_BIT_OFFSET = 0;
  localparam int STATIC_REG1_RD_ALLOW_FULL_BURST_BIT_WIDTH = 1;
  localparam bit STATIC_REG1_RD_ALLOW_FULL_BURST_BIT_MASK = 1'h1;
  localparam int STATIC_REG1_RD_ALLOW_FULL_BURST_BIT_OFFSET = 12;
  localparam int STATIC_REG1_RD_ALLOW_FULL_FIFO_BIT_WIDTH = 1;
  localparam bit STATIC_REG1_RD_ALLOW_FULL_FIFO_BIT_MASK = 1'h1;
  localparam int STATIC_REG1_RD_ALLOW_FULL_FIFO_BIT_OFFSET = 13;
  localparam int STATIC_REG1_RD_TOKENS_BIT_WIDTH = 6;
  localparam bit [5:0] STATIC_REG1_RD_TOKENS_BIT_MASK = 6'h3f;
  localparam int STATIC_REG1_RD_TOKENS_BIT_OFFSET = 16;
  localparam int STATIC_REG1_RD_OUTS_MAX_BIT_WIDTH = 4;
  localparam bit [3:0] STATIC_REG1_RD_OUTS_MAX_BIT_MASK = 4'hf;
  localparam int STATIC_REG1_RD_OUTS_MAX_BIT_OFFSET = 24;
  localparam int STATIC_REG1_RD_OUTSTANDING_BIT_WIDTH = 1;
  localparam bit STATIC_REG1_RD_OUTSTANDING_BIT_MASK = 1'h1;
  localparam int STATIC_REG1_RD_OUTSTANDING_BIT_OFFSET = 30;
  localparam int STATIC_REG1_RD_INCR_BIT_WIDTH = 1;
  localparam bit STATIC_REG1_RD_INCR_BIT_MASK = 1'h1;
  localparam int STATIC_REG1_RD_INCR_BIT_OFFSET = 31;
  localparam int STATIC_REG2_BYTE_WIDTH = 4;
  localparam int STATIC_REG2_BYTE_SIZE = 4;
  localparam bit [12:0] STATIC_REG2_BYTE_OFFSET = 13'h0018;
  localparam int STATIC_REG2_FRAME_WIDTH_BIT_WIDTH = 12;
  localparam bit [11:0] STATIC_REG2_FRAME_WIDTH_BIT_MASK = 12'hfff;
  localparam int STATIC_REG2_FRAME_WIDTH_BIT_OFFSET = 0;
  localparam int STATIC_REG2_BLOCK_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_BLOCK_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_BLOCK_BIT_OFFSET = 15;
  localparam int STATIC_REG2_JOINT_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_JOINT_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_JOINT_BIT_OFFSET = 16;
  localparam int STATIC_REG2_AUTO_RETRY_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_AUTO_RETRY_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_AUTO_RETRY_BIT_OFFSET = 17;
  localparam int STATIC_REG2_RD_CMD_PORT_NUM_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_RD_CMD_PORT_NUM_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_RD_CMD_PORT_NUM_BIT_OFFSET = 20;
  localparam int STATIC_REG2_RD_PORT_NUM_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_RD_PORT_NUM_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_RD_PORT_NUM_BIT_OFFSET = 21;
  localparam int STATIC_REG2_WR_PORT_NUM_BIT_WIDTH = 1;
  localparam bit STATIC_REG2_WR_PORT_NUM_BIT_MASK = 1'h1;
  localparam int STATIC_REG2_WR_PORT_NUM_BIT_OFFSET = 22;
  localparam int STATIC_REG2_INT_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] STATIC_REG2_INT_NUM_BIT_MASK = 3'h7;
  localparam int STATIC_REG2_INT_NUM_BIT_OFFSET = 24;
  localparam int STATIC_REG2_END_SWAP_BIT_WIDTH = 2;
  localparam bit [1:0] STATIC_REG2_END_SWAP_BIT_MASK = 2'h3;
  localparam int STATIC_REG2_END_SWAP_BIT_OFFSET = 28;
  localparam int STATIC_REG3_BYTE_WIDTH = 4;
  localparam int STATIC_REG3_BYTE_SIZE = 4;
  localparam bit [12:0] STATIC_REG3_BYTE_OFFSET = 13'h001c;
  localparam int STATIC_REG3_RD_WAIT_LIMIT_BIT_WIDTH = 12;
  localparam bit [11:0] STATIC_REG3_RD_WAIT_LIMIT_BIT_MASK = 12'hfff;
  localparam int STATIC_REG3_RD_WAIT_LIMIT_BIT_OFFSET = 0;
  localparam int STATIC_REG3_WR_WAIT_LIMIT_BIT_WIDTH = 12;
  localparam bit [11:0] STATIC_REG3_WR_WAIT_LIMIT_BIT_MASK = 12'hfff;
  localparam int STATIC_REG3_WR_WAIT_LIMIT_BIT_OFFSET = 16;
  localparam int STATIC_REG4_BYTE_WIDTH = 4;
  localparam int STATIC_REG4_BYTE_SIZE = 4;
  localparam bit [12:0] STATIC_REG4_BYTE_OFFSET = 13'h0020;
  localparam int STATIC_REG4_RD_PERIPH_NUM_BIT_WIDTH = 5;
  localparam bit [4:0] STATIC_REG4_RD_PERIPH_NUM_BIT_MASK = 5'h1f;
  localparam int STATIC_REG4_RD_PERIPH_NUM_BIT_OFFSET = 0;
  localparam int STATIC_REG4_RD_PERIPH_DELAY_BIT_WIDTH = 3;
  localparam bit [2:0] STATIC_REG4_RD_PERIPH_DELAY_BIT_MASK = 3'h7;
  localparam int STATIC_REG4_RD_PERIPH_DELAY_BIT_OFFSET = 8;
  localparam int STATIC_REG4_RD_PERIPH_BLOCK_BIT_WIDTH = 1;
  localparam bit STATIC_REG4_RD_PERIPH_BLOCK_BIT_MASK = 1'h1;
  localparam int STATIC_REG4_RD_PERIPH_BLOCK_BIT_OFFSET = 15;
  localparam int STATIC_REG4_WR_PERIPH_NUM_BIT_WIDTH = 5;
  localparam bit [4:0] STATIC_REG4_WR_PERIPH_NUM_BIT_MASK = 5'h1f;
  localparam int STATIC_REG4_WR_PERIPH_NUM_BIT_OFFSET = 16;
  localparam int STATIC_REG4_WR_PERIPH_DELAY_BIT_WIDTH = 3;
  localparam bit [2:0] STATIC_REG4_WR_PERIPH_DELAY_BIT_MASK = 3'h7;
  localparam int STATIC_REG4_WR_PERIPH_DELAY_BIT_OFFSET = 24;
  localparam int STATIC_REG4_WR_PERIPH_BLOCK_BIT_WIDTH = 1;
  localparam bit STATIC_REG4_WR_PERIPH_BLOCK_BIT_MASK = 1'h1;
  localparam int STATIC_REG4_WR_PERIPH_BLOCK_BIT_OFFSET = 31;
  localparam int RESTRICT_REG_BYTE_WIDTH = 4;
  localparam int RESTRICT_REG_BYTE_SIZE = 4;
  localparam bit [12:0] RESTRICT_REG_BYTE_OFFSET = 13'h002c;
  localparam int RESTRICT_REG_RD_ALLOW_FULL_FIFO_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_RD_ALLOW_FULL_FIFO_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_RD_ALLOW_FULL_FIFO_BIT_OFFSET = 0;
  localparam int RESTRICT_REG_WR_ALLOW_FULL_FIFO_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_WR_ALLOW_FULL_FIFO_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_WR_ALLOW_FULL_FIFO_BIT_OFFSET = 1;
  localparam int RESTRICT_REG_ALLOW_FULL_FIFO_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_ALLOW_FULL_FIFO_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_ALLOW_FULL_FIFO_BIT_OFFSET = 2;
  localparam int RESTRICT_REG_ALLOW_FULL_BURST_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_ALLOW_FULL_BURST_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_ALLOW_FULL_BURST_BIT_OFFSET = 3;
  localparam int RESTRICT_REG_ALLOW_JOINT_BURST_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_ALLOW_JOINT_BURST_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_ALLOW_JOINT_BURST_BIT_OFFSET = 4;
  localparam int RESTRICT_REG_RD_OUTSTANDING_STAT_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_RD_OUTSTANDING_STAT_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_RD_OUTSTANDING_STAT_BIT_OFFSET = 5;
  localparam int RESTRICT_REG_WR_OUTSTANDING_STAT_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_WR_OUTSTANDING_STAT_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_WR_OUTSTANDING_STAT_BIT_OFFSET = 6;
  localparam int RESTRICT_REG_BLOCK_NON_ALIGN_STAT_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_BLOCK_NON_ALIGN_STAT_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_BLOCK_NON_ALIGN_STAT_BIT_OFFSET = 7;
  localparam int RESTRICT_REG_SIMPLE_STAT_BIT_WIDTH = 1;
  localparam bit RESTRICT_REG_SIMPLE_STAT_BIT_MASK = 1'h1;
  localparam int RESTRICT_REG_SIMPLE_STAT_BIT_OFFSET = 8;
  localparam int READ_OFFSET_REG_BYTE_WIDTH = 4;
  localparam int READ_OFFSET_REG_BYTE_SIZE = 4;
  localparam bit [12:0] READ_OFFSET_REG_BYTE_OFFSET = 13'h0030;
  localparam int READ_OFFSET_REG_RD_OFFSET_BIT_WIDTH = 16;
  localparam bit [15:0] READ_OFFSET_REG_RD_OFFSET_BIT_MASK = 16'hffff;
  localparam int READ_OFFSET_REG_RD_OFFSET_BIT_OFFSET = 0;
  localparam int WRITE_OFFSET_REG_BYTE_WIDTH = 4;
  localparam int WRITE_OFFSET_REG_BYTE_SIZE = 4;
  localparam bit [12:0] WRITE_OFFSET_REG_BYTE_OFFSET = 13'h0034;
  localparam int WRITE_OFFSET_REG_WR_OFFSET_BIT_WIDTH = 16;
  localparam bit [15:0] WRITE_OFFSET_REG_WR_OFFSET_BIT_MASK = 16'hffff;
  localparam int WRITE_OFFSET_REG_WR_OFFSET_BIT_OFFSET = 0;
  localparam int FIFO_FULLNESS_REG_BYTE_WIDTH = 4;
  localparam int FIFO_FULLNESS_REG_BYTE_SIZE = 4;
  localparam bit [12:0] FIFO_FULLNESS_REG_BYTE_OFFSET = 13'h0038;
  localparam int FIFO_FULLNESS_REG_RD_GAP_BIT_WIDTH = 10;
  localparam bit [9:0] FIFO_FULLNESS_REG_RD_GAP_BIT_MASK = 10'h3ff;
  localparam int FIFO_FULLNESS_REG_RD_GAP_BIT_OFFSET = 0;
  localparam int FIFO_FULLNESS_REG_WR_FULLNESS_BIT_WIDTH = 10;
  localparam bit [9:0] FIFO_FULLNESS_REG_WR_FULLNESS_BIT_MASK = 10'h3ff;
  localparam int FIFO_FULLNESS_REG_WR_FULLNESS_BIT_OFFSET = 16;
  localparam int CMD_OUTS_REG_BYTE_WIDTH = 4;
  localparam int CMD_OUTS_REG_BYTE_SIZE = 4;
  localparam bit [12:0] CMD_OUTS_REG_BYTE_OFFSET = 13'h003c;
  localparam int CMD_OUTS_REG_RD_CMD_OUTS_BIT_WIDTH = 6;
  localparam bit [5:0] CMD_OUTS_REG_RD_CMD_OUTS_BIT_MASK = 6'h3f;
  localparam int CMD_OUTS_REG_RD_CMD_OUTS_BIT_OFFSET = 0;
  localparam int CMD_OUTS_REG_WR_CMD_OUTS_BIT_WIDTH = 6;
  localparam bit [5:0] CMD_OUTS_REG_WR_CMD_OUTS_BIT_MASK = 6'h3f;
  localparam int CMD_OUTS_REG_WR_CMD_OUTS_BIT_OFFSET = 8;
  localparam int CH_ENABLE_REG_BYTE_WIDTH = 4;
  localparam int CH_ENABLE_REG_BYTE_SIZE = 4;
  localparam bit [12:0] CH_ENABLE_REG_BYTE_OFFSET = 13'h0040;
  localparam int CH_ENABLE_REG_CH_ENABLE_BIT_WIDTH = 1;
  localparam bit CH_ENABLE_REG_CH_ENABLE_BIT_MASK = 1'h1;
  localparam int CH_ENABLE_REG_CH_ENABLE_BIT_OFFSET = 0;
  localparam int CH_START_REG_BYTE_WIDTH = 4;
  localparam int CH_START_REG_BYTE_SIZE = 4;
  localparam bit [12:0] CH_START_REG_BYTE_OFFSET = 13'h0044;
  localparam int CH_START_REG_CH_START_BIT_WIDTH = 1;
  localparam bit CH_START_REG_CH_START_BIT_MASK = 1'h1;
  localparam int CH_START_REG_CH_START_BIT_OFFSET = 0;
  localparam int CH_ACTIVE_REG_BYTE_WIDTH = 4;
  localparam int CH_ACTIVE_REG_BYTE_SIZE = 4;
  localparam bit [12:0] CH_ACTIVE_REG_BYTE_OFFSET = 13'h0048;
  localparam int CH_ACTIVE_REG_CH_RD_ACTIVE_BIT_WIDTH = 1;
  localparam bit CH_ACTIVE_REG_CH_RD_ACTIVE_BIT_MASK = 1'h1;
  localparam int CH_ACTIVE_REG_CH_RD_ACTIVE_BIT_OFFSET = 0;
  localparam int CH_ACTIVE_REG_CH_WR_ACTIVE_BIT_WIDTH = 1;
  localparam bit CH_ACTIVE_REG_CH_WR_ACTIVE_BIT_MASK = 1'h1;
  localparam int CH_ACTIVE_REG_CH_WR_ACTIVE_BIT_OFFSET = 1;
  localparam int COUNT_REG_BYTE_WIDTH = 4;
  localparam int COUNT_REG_BYTE_SIZE = 4;
  localparam bit [12:0] COUNT_REG_BYTE_OFFSET = 13'h0050;
  localparam int COUNT_REG_BUFF_COUNT_BIT_WIDTH = 16;
  localparam bit [15:0] COUNT_REG_BUFF_COUNT_BIT_MASK = 16'hffff;
  localparam int COUNT_REG_BUFF_COUNT_BIT_OFFSET = 0;
  localparam int COUNT_REG_INT_COUNT_BIT_WIDTH = 6;
  localparam bit [5:0] COUNT_REG_INT_COUNT_BIT_MASK = 6'h3f;
  localparam int COUNT_REG_INT_COUNT_BIT_OFFSET = 16;
  localparam int INT_RAWSTAT_REG_BYTE_WIDTH = 4;
  localparam int INT_RAWSTAT_REG_BYTE_SIZE = 4;
  localparam bit [12:0] INT_RAWSTAT_REG_BYTE_OFFSET = 13'h00a0;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_CH_END_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_CH_END_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_CH_END_BIT_OFFSET = 0;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_RD_DECERR_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_RD_DECERR_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_RD_DECERR_BIT_OFFSET = 1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_RD_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_RD_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_RD_SLVERR_BIT_OFFSET = 2;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WR_DECERR_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_WR_DECERR_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WR_DECERR_BIT_OFFSET = 3;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WR_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_WR_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WR_SLVERR_BIT_OFFSET = 4;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_OVERFLOW_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_OVERFLOW_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_OVERFLOW_BIT_OFFSET = 5;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_UNDERFLOW_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_UNDERFLOW_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_UNDERFLOW_BIT_OFFSET = 6;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_R_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_R_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_R_BIT_OFFSET = 7;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AR_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AR_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AR_BIT_OFFSET = 8;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_B_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_B_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_B_BIT_OFFSET = 9;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_W_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_W_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_W_BIT_OFFSET = 10;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AW_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AW_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_TIMEOUT_AW_BIT_OFFSET = 11;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WDT_BIT_WIDTH = 1;
  localparam bit INT_RAWSTAT_REG_INT_RAWSTAT_WDT_BIT_MASK = 1'h1;
  localparam int INT_RAWSTAT_REG_INT_RAWSTAT_WDT_BIT_OFFSET = 12;
  localparam int INT_CLEAR_REG_BYTE_WIDTH = 4;
  localparam int INT_CLEAR_REG_BYTE_SIZE = 4;
  localparam bit [12:0] INT_CLEAR_REG_BYTE_OFFSET = 13'h00a4;
  localparam int INT_CLEAR_REG_INT_CLR_CH_END_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_CH_END_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_CH_END_BIT_OFFSET = 0;
  localparam int INT_CLEAR_REG_INT_CLR_RD_DECERR_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_RD_DECERR_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_RD_DECERR_BIT_OFFSET = 1;
  localparam int INT_CLEAR_REG_INT_CLR_RD_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_RD_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_RD_SLVERR_BIT_OFFSET = 2;
  localparam int INT_CLEAR_REG_INT_CLR_WR_DECERR_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_WR_DECERR_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_WR_DECERR_BIT_OFFSET = 3;
  localparam int INT_CLEAR_REG_INT_CLR_WR_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_WR_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_WR_SLVERR_BIT_OFFSET = 4;
  localparam int INT_CLEAR_REG_INT_CLR_OVERFLOW_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_OVERFLOW_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_OVERFLOW_BIT_OFFSET = 5;
  localparam int INT_CLEAR_REG_INT_CLR_UNDERFLOW_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_UNDERFLOW_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_UNDERFLOW_BIT_OFFSET = 6;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_R_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_TIMEOUT_R_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_R_BIT_OFFSET = 7;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_AR_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_TIMEOUT_AR_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_AR_BIT_OFFSET = 8;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_B_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_TIMEOUT_B_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_B_BIT_OFFSET = 9;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_W_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_TIMEOUT_W_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_W_BIT_OFFSET = 10;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_AW_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_TIMEOUT_AW_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_TIMEOUT_AW_BIT_OFFSET = 11;
  localparam int INT_CLEAR_REG_INT_CLR_WDT_BIT_WIDTH = 1;
  localparam bit INT_CLEAR_REG_INT_CLR_WDT_BIT_MASK = 1'h1;
  localparam int INT_CLEAR_REG_INT_CLR_WDT_BIT_OFFSET = 12;
  localparam int INT_ENABLE_REG_BYTE_WIDTH = 4;
  localparam int INT_ENABLE_REG_BYTE_SIZE = 4;
  localparam bit [12:0] INT_ENABLE_REG_BYTE_OFFSET = 13'h00a8;
  localparam int INT_ENABLE_REG_INT_ENABLE_CH_END_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_CH_END_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_CH_END_BIT_OFFSET = 0;
  localparam int INT_ENABLE_REG_INT_ENABLE_RD_DECERR_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_RD_DECERR_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_RD_DECERR_BIT_OFFSET = 1;
  localparam int INT_ENABLE_REG_INT_ENABLE_RD_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_RD_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_RD_SLVERR_BIT_OFFSET = 2;
  localparam int INT_ENABLE_REG_INT_ENABLE_WR_DECERR_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_WR_DECERR_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_WR_DECERR_BIT_OFFSET = 3;
  localparam int INT_ENABLE_REG_INT_ENABLE_WR_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_WR_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_WR_SLVERR_BIT_OFFSET = 4;
  localparam int INT_ENABLE_REG_INT_ENABLE_OVERFLOW_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_OVERFLOW_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_OVERFLOW_BIT_OFFSET = 5;
  localparam int INT_ENABLE_REG_INT_ENABLE_UNDERFLOW_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_UNDERFLOW_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_UNDERFLOW_BIT_OFFSET = 6;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_R_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_TIMEOUT_R_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_R_BIT_OFFSET = 7;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AR_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AR_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AR_BIT_OFFSET = 8;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_B_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_TIMEOUT_B_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_B_BIT_OFFSET = 9;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_W_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_TIMEOUT_W_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_W_BIT_OFFSET = 10;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AW_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AW_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_TIMEOUT_AW_BIT_OFFSET = 11;
  localparam int INT_ENABLE_REG_INT_ENABLE_WDT_BIT_WIDTH = 1;
  localparam bit INT_ENABLE_REG_INT_ENABLE_WDT_BIT_MASK = 1'h1;
  localparam int INT_ENABLE_REG_INT_ENABLE_WDT_BIT_OFFSET = 12;
  localparam int INT_STATUS_REG_BYTE_WIDTH = 4;
  localparam int INT_STATUS_REG_BYTE_SIZE = 4;
  localparam bit [12:0] INT_STATUS_REG_BYTE_OFFSET = 13'h00ac;
  localparam int INT_STATUS_REG_INT_STATUS_CH_END_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_CH_END_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_CH_END_BIT_OFFSET = 0;
  localparam int INT_STATUS_REG_INT_STATUS_RD_DECERR_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_RD_DECERR_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_RD_DECERR_BIT_OFFSET = 1;
  localparam int INT_STATUS_REG_INT_STATUS_RD_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_RD_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_RD_SLVERR_BIT_OFFSET = 2;
  localparam int INT_STATUS_REG_INT_STATUS_WR_DECERR_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_WR_DECERR_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_WR_DECERR_BIT_OFFSET = 3;
  localparam int INT_STATUS_REG_INT_STATUS_WR_SLVERR_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_WR_SLVERR_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_WR_SLVERR_BIT_OFFSET = 4;
  localparam int INT_STATUS_REG_INT_STATUS_OVERFLOW_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_OVERFLOW_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_OVERFLOW_BIT_OFFSET = 5;
  localparam int INT_STATUS_REG_INT_STATUS_UNDERFLOW_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_UNDERFLOW_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_UNDERFLOW_BIT_OFFSET = 6;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_R_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_TIMEOUT_R_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_R_BIT_OFFSET = 7;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_AR_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_TIMEOUT_AR_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_AR_BIT_OFFSET = 8;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_B_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_TIMEOUT_B_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_B_BIT_OFFSET = 9;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_W_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_TIMEOUT_W_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_W_BIT_OFFSET = 10;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_AW_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_TIMEOUT_AW_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_TIMEOUT_AW_BIT_OFFSET = 11;
  localparam int INT_STATUS_REG_INT_STATUS_WDT_BIT_WIDTH = 1;
  localparam bit INT_STATUS_REG_INT_STATUS_WDT_BIT_MASK = 1'h1;
  localparam int INT_STATUS_REG_INT_STATUS_WDT_BIT_OFFSET = 12;
  localparam int INT0_STATUS_BYTE_WIDTH = 4;
  localparam int INT0_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT0_STATUS_BYTE_OFFSET = 13'h1000;
  localparam int INT0_STATUS_CORE0_CH0_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH0_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH0_INT0_STAT_BIT_OFFSET = 0;
  localparam int INT0_STATUS_CORE0_CH1_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH1_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH1_INT0_STAT_BIT_OFFSET = 1;
  localparam int INT0_STATUS_CORE0_CH2_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH2_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH2_INT0_STAT_BIT_OFFSET = 2;
  localparam int INT0_STATUS_CORE0_CH3_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH3_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH3_INT0_STAT_BIT_OFFSET = 3;
  localparam int INT0_STATUS_CORE0_CH4_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH4_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH4_INT0_STAT_BIT_OFFSET = 4;
  localparam int INT0_STATUS_CORE0_CH5_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH5_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH5_INT0_STAT_BIT_OFFSET = 5;
  localparam int INT0_STATUS_CORE0_CH6_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH6_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH6_INT0_STAT_BIT_OFFSET = 6;
  localparam int INT0_STATUS_CORE0_CH7_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE0_CH7_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE0_CH7_INT0_STAT_BIT_OFFSET = 7;
  localparam int INT0_STATUS_CORE1_CH0_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH0_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH0_INT0_STAT_BIT_OFFSET = 8;
  localparam int INT0_STATUS_CORE1_CH1_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH1_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH1_INT0_STAT_BIT_OFFSET = 9;
  localparam int INT0_STATUS_CORE1_CH2_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH2_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH2_INT0_STAT_BIT_OFFSET = 10;
  localparam int INT0_STATUS_CORE1_CH3_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH3_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH3_INT0_STAT_BIT_OFFSET = 11;
  localparam int INT0_STATUS_CORE1_CH4_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH4_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH4_INT0_STAT_BIT_OFFSET = 12;
  localparam int INT0_STATUS_CORE1_CH5_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH5_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH5_INT0_STAT_BIT_OFFSET = 13;
  localparam int INT0_STATUS_CORE1_CH6_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH6_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH6_INT0_STAT_BIT_OFFSET = 14;
  localparam int INT0_STATUS_CORE1_CH7_INT0_STAT_BIT_WIDTH = 1;
  localparam bit INT0_STATUS_CORE1_CH7_INT0_STAT_BIT_MASK = 1'h1;
  localparam int INT0_STATUS_CORE1_CH7_INT0_STAT_BIT_OFFSET = 15;
  localparam int INT1_STATUS_BYTE_WIDTH = 4;
  localparam int INT1_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT1_STATUS_BYTE_OFFSET = 13'h1004;
  localparam int INT1_STATUS_CORE0_CH0_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH0_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH0_INT1_STAT_BIT_OFFSET = 0;
  localparam int INT1_STATUS_CORE0_CH1_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH1_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH1_INT1_STAT_BIT_OFFSET = 1;
  localparam int INT1_STATUS_CORE0_CH2_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH2_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH2_INT1_STAT_BIT_OFFSET = 2;
  localparam int INT1_STATUS_CORE0_CH3_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH3_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH3_INT1_STAT_BIT_OFFSET = 3;
  localparam int INT1_STATUS_CORE0_CH4_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH4_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH4_INT1_STAT_BIT_OFFSET = 4;
  localparam int INT1_STATUS_CORE0_CH5_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH5_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH5_INT1_STAT_BIT_OFFSET = 5;
  localparam int INT1_STATUS_CORE0_CH6_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH6_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH6_INT1_STAT_BIT_OFFSET = 6;
  localparam int INT1_STATUS_CORE0_CH7_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE0_CH7_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE0_CH7_INT1_STAT_BIT_OFFSET = 7;
  localparam int INT1_STATUS_CORE1_CH0_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH0_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH0_INT1_STAT_BIT_OFFSET = 8;
  localparam int INT1_STATUS_CORE1_CH1_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH1_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH1_INT1_STAT_BIT_OFFSET = 9;
  localparam int INT1_STATUS_CORE1_CH2_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH2_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH2_INT1_STAT_BIT_OFFSET = 10;
  localparam int INT1_STATUS_CORE1_CH3_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH3_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH3_INT1_STAT_BIT_OFFSET = 11;
  localparam int INT1_STATUS_CORE1_CH4_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH4_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH4_INT1_STAT_BIT_OFFSET = 12;
  localparam int INT1_STATUS_CORE1_CH5_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH5_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH5_INT1_STAT_BIT_OFFSET = 13;
  localparam int INT1_STATUS_CORE1_CH6_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH6_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH6_INT1_STAT_BIT_OFFSET = 14;
  localparam int INT1_STATUS_CORE1_CH7_INT1_STAT_BIT_WIDTH = 1;
  localparam bit INT1_STATUS_CORE1_CH7_INT1_STAT_BIT_MASK = 1'h1;
  localparam int INT1_STATUS_CORE1_CH7_INT1_STAT_BIT_OFFSET = 15;
  localparam int INT2_STATUS_BYTE_WIDTH = 4;
  localparam int INT2_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT2_STATUS_BYTE_OFFSET = 13'h1008;
  localparam int INT2_STATUS_CORE0_CH0_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH0_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH0_INT2_STAT_BIT_OFFSET = 0;
  localparam int INT2_STATUS_CORE0_CH1_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH1_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH1_INT2_STAT_BIT_OFFSET = 1;
  localparam int INT2_STATUS_CORE0_CH2_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH2_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH2_INT2_STAT_BIT_OFFSET = 2;
  localparam int INT2_STATUS_CORE0_CH3_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH3_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH3_INT2_STAT_BIT_OFFSET = 3;
  localparam int INT2_STATUS_CORE0_CH4_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH4_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH4_INT2_STAT_BIT_OFFSET = 4;
  localparam int INT2_STATUS_CORE0_CH5_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH5_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH5_INT2_STAT_BIT_OFFSET = 5;
  localparam int INT2_STATUS_CORE0_CH6_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH6_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH6_INT2_STAT_BIT_OFFSET = 6;
  localparam int INT2_STATUS_CORE0_CH7_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE0_CH7_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE0_CH7_INT2_STAT_BIT_OFFSET = 7;
  localparam int INT2_STATUS_CORE1_CH0_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH0_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH0_INT2_STAT_BIT_OFFSET = 8;
  localparam int INT2_STATUS_CORE1_CH1_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH1_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH1_INT2_STAT_BIT_OFFSET = 9;
  localparam int INT2_STATUS_CORE1_CH2_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH2_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH2_INT2_STAT_BIT_OFFSET = 10;
  localparam int INT2_STATUS_CORE1_CH3_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH3_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH3_INT2_STAT_BIT_OFFSET = 11;
  localparam int INT2_STATUS_CORE1_CH4_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH4_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH4_INT2_STAT_BIT_OFFSET = 12;
  localparam int INT2_STATUS_CORE1_CH5_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH5_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH5_INT2_STAT_BIT_OFFSET = 13;
  localparam int INT2_STATUS_CORE1_CH6_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH6_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH6_INT2_STAT_BIT_OFFSET = 14;
  localparam int INT2_STATUS_CORE1_CH7_INT2_STAT_BIT_WIDTH = 1;
  localparam bit INT2_STATUS_CORE1_CH7_INT2_STAT_BIT_MASK = 1'h1;
  localparam int INT2_STATUS_CORE1_CH7_INT2_STAT_BIT_OFFSET = 15;
  localparam int INT3_STATUS_BYTE_WIDTH = 4;
  localparam int INT3_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT3_STATUS_BYTE_OFFSET = 13'h100c;
  localparam int INT3_STATUS_CORE0_CH0_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH0_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH0_INT3_STAT_BIT_OFFSET = 0;
  localparam int INT3_STATUS_CORE0_CH1_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH1_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH1_INT3_STAT_BIT_OFFSET = 1;
  localparam int INT3_STATUS_CORE0_CH2_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH2_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH2_INT3_STAT_BIT_OFFSET = 2;
  localparam int INT3_STATUS_CORE0_CH3_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH3_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH3_INT3_STAT_BIT_OFFSET = 3;
  localparam int INT3_STATUS_CORE0_CH4_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH4_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH4_INT3_STAT_BIT_OFFSET = 4;
  localparam int INT3_STATUS_CORE0_CH5_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH5_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH5_INT3_STAT_BIT_OFFSET = 5;
  localparam int INT3_STATUS_CORE0_CH6_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH6_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH6_INT3_STAT_BIT_OFFSET = 6;
  localparam int INT3_STATUS_CORE0_CH7_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE0_CH7_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE0_CH7_INT3_STAT_BIT_OFFSET = 7;
  localparam int INT3_STATUS_CORE1_CH0_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH0_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH0_INT3_STAT_BIT_OFFSET = 8;
  localparam int INT3_STATUS_CORE1_CH1_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH1_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH1_INT3_STAT_BIT_OFFSET = 9;
  localparam int INT3_STATUS_CORE1_CH2_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH2_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH2_INT3_STAT_BIT_OFFSET = 10;
  localparam int INT3_STATUS_CORE1_CH3_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH3_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH3_INT3_STAT_BIT_OFFSET = 11;
  localparam int INT3_STATUS_CORE1_CH4_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH4_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH4_INT3_STAT_BIT_OFFSET = 12;
  localparam int INT3_STATUS_CORE1_CH5_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH5_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH5_INT3_STAT_BIT_OFFSET = 13;
  localparam int INT3_STATUS_CORE1_CH6_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH6_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH6_INT3_STAT_BIT_OFFSET = 14;
  localparam int INT3_STATUS_CORE1_CH7_INT3_STAT_BIT_WIDTH = 1;
  localparam bit INT3_STATUS_CORE1_CH7_INT3_STAT_BIT_MASK = 1'h1;
  localparam int INT3_STATUS_CORE1_CH7_INT3_STAT_BIT_OFFSET = 15;
  localparam int INT4_STATUS_BYTE_WIDTH = 4;
  localparam int INT4_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT4_STATUS_BYTE_OFFSET = 13'h1010;
  localparam int INT4_STATUS_CORE0_CH0_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH0_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH0_INT4_STAT_BIT_OFFSET = 0;
  localparam int INT4_STATUS_CORE0_CH1_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH1_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH1_INT4_STAT_BIT_OFFSET = 1;
  localparam int INT4_STATUS_CORE0_CH2_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH2_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH2_INT4_STAT_BIT_OFFSET = 2;
  localparam int INT4_STATUS_CORE0_CH3_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH3_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH3_INT4_STAT_BIT_OFFSET = 3;
  localparam int INT4_STATUS_CORE0_CH4_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH4_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH4_INT4_STAT_BIT_OFFSET = 4;
  localparam int INT4_STATUS_CORE0_CH5_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH5_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH5_INT4_STAT_BIT_OFFSET = 5;
  localparam int INT4_STATUS_CORE0_CH6_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH6_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH6_INT4_STAT_BIT_OFFSET = 6;
  localparam int INT4_STATUS_CORE0_CH7_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE0_CH7_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE0_CH7_INT4_STAT_BIT_OFFSET = 7;
  localparam int INT4_STATUS_CORE1_CH0_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH0_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH0_INT4_STAT_BIT_OFFSET = 8;
  localparam int INT4_STATUS_CORE1_CH1_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH1_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH1_INT4_STAT_BIT_OFFSET = 9;
  localparam int INT4_STATUS_CORE1_CH2_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH2_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH2_INT4_STAT_BIT_OFFSET = 10;
  localparam int INT4_STATUS_CORE1_CH3_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH3_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH3_INT4_STAT_BIT_OFFSET = 11;
  localparam int INT4_STATUS_CORE1_CH4_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH4_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH4_INT4_STAT_BIT_OFFSET = 12;
  localparam int INT4_STATUS_CORE1_CH5_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH5_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH5_INT4_STAT_BIT_OFFSET = 13;
  localparam int INT4_STATUS_CORE1_CH6_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH6_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH6_INT4_STAT_BIT_OFFSET = 14;
  localparam int INT4_STATUS_CORE1_CH7_INT4_STAT_BIT_WIDTH = 1;
  localparam bit INT4_STATUS_CORE1_CH7_INT4_STAT_BIT_MASK = 1'h1;
  localparam int INT4_STATUS_CORE1_CH7_INT4_STAT_BIT_OFFSET = 15;
  localparam int INT5_STATUS_BYTE_WIDTH = 4;
  localparam int INT5_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT5_STATUS_BYTE_OFFSET = 13'h1014;
  localparam int INT5_STATUS_CORE0_CH0_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH0_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH0_INT5_STAT_BIT_OFFSET = 0;
  localparam int INT5_STATUS_CORE0_CH1_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH1_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH1_INT5_STAT_BIT_OFFSET = 1;
  localparam int INT5_STATUS_CORE0_CH2_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH2_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH2_INT5_STAT_BIT_OFFSET = 2;
  localparam int INT5_STATUS_CORE0_CH3_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH3_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH3_INT5_STAT_BIT_OFFSET = 3;
  localparam int INT5_STATUS_CORE0_CH4_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH4_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH4_INT5_STAT_BIT_OFFSET = 4;
  localparam int INT5_STATUS_CORE0_CH5_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH5_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH5_INT5_STAT_BIT_OFFSET = 5;
  localparam int INT5_STATUS_CORE0_CH6_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH6_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH6_INT5_STAT_BIT_OFFSET = 6;
  localparam int INT5_STATUS_CORE0_CH7_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE0_CH7_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE0_CH7_INT5_STAT_BIT_OFFSET = 7;
  localparam int INT5_STATUS_CORE1_CH0_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH0_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH0_INT5_STAT_BIT_OFFSET = 8;
  localparam int INT5_STATUS_CORE1_CH1_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH1_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH1_INT5_STAT_BIT_OFFSET = 9;
  localparam int INT5_STATUS_CORE1_CH2_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH2_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH2_INT5_STAT_BIT_OFFSET = 10;
  localparam int INT5_STATUS_CORE1_CH3_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH3_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH3_INT5_STAT_BIT_OFFSET = 11;
  localparam int INT5_STATUS_CORE1_CH4_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH4_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH4_INT5_STAT_BIT_OFFSET = 12;
  localparam int INT5_STATUS_CORE1_CH5_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH5_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH5_INT5_STAT_BIT_OFFSET = 13;
  localparam int INT5_STATUS_CORE1_CH6_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH6_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH6_INT5_STAT_BIT_OFFSET = 14;
  localparam int INT5_STATUS_CORE1_CH7_INT5_STAT_BIT_WIDTH = 1;
  localparam bit INT5_STATUS_CORE1_CH7_INT5_STAT_BIT_MASK = 1'h1;
  localparam int INT5_STATUS_CORE1_CH7_INT5_STAT_BIT_OFFSET = 15;
  localparam int INT6_STATUS_BYTE_WIDTH = 4;
  localparam int INT6_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT6_STATUS_BYTE_OFFSET = 13'h1018;
  localparam int INT6_STATUS_CORE0_CH0_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH0_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH0_INT6_STAT_BIT_OFFSET = 0;
  localparam int INT6_STATUS_CORE0_CH1_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH1_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH1_INT6_STAT_BIT_OFFSET = 1;
  localparam int INT6_STATUS_CORE0_CH2_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH2_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH2_INT6_STAT_BIT_OFFSET = 2;
  localparam int INT6_STATUS_CORE0_CH3_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH3_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH3_INT6_STAT_BIT_OFFSET = 3;
  localparam int INT6_STATUS_CORE0_CH4_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH4_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH4_INT6_STAT_BIT_OFFSET = 4;
  localparam int INT6_STATUS_CORE0_CH5_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH5_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH5_INT6_STAT_BIT_OFFSET = 5;
  localparam int INT6_STATUS_CORE0_CH6_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH6_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH6_INT6_STAT_BIT_OFFSET = 6;
  localparam int INT6_STATUS_CORE0_CH7_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE0_CH7_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE0_CH7_INT6_STAT_BIT_OFFSET = 7;
  localparam int INT6_STATUS_CORE1_CH0_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH0_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH0_INT6_STAT_BIT_OFFSET = 8;
  localparam int INT6_STATUS_CORE1_CH1_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH1_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH1_INT6_STAT_BIT_OFFSET = 9;
  localparam int INT6_STATUS_CORE1_CH2_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH2_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH2_INT6_STAT_BIT_OFFSET = 10;
  localparam int INT6_STATUS_CORE1_CH3_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH3_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH3_INT6_STAT_BIT_OFFSET = 11;
  localparam int INT6_STATUS_CORE1_CH4_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH4_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH4_INT6_STAT_BIT_OFFSET = 12;
  localparam int INT6_STATUS_CORE1_CH5_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH5_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH5_INT6_STAT_BIT_OFFSET = 13;
  localparam int INT6_STATUS_CORE1_CH6_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH6_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH6_INT6_STAT_BIT_OFFSET = 14;
  localparam int INT6_STATUS_CORE1_CH7_INT6_STAT_BIT_WIDTH = 1;
  localparam bit INT6_STATUS_CORE1_CH7_INT6_STAT_BIT_MASK = 1'h1;
  localparam int INT6_STATUS_CORE1_CH7_INT6_STAT_BIT_OFFSET = 15;
  localparam int INT7_STATUS_BYTE_WIDTH = 4;
  localparam int INT7_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] INT7_STATUS_BYTE_OFFSET = 13'h101c;
  localparam int INT7_STATUS_CORE0_CH0_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH0_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH0_INT7_STAT_BIT_OFFSET = 0;
  localparam int INT7_STATUS_CORE0_CH1_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH1_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH1_INT7_STAT_BIT_OFFSET = 1;
  localparam int INT7_STATUS_CORE0_CH2_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH2_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH2_INT7_STAT_BIT_OFFSET = 2;
  localparam int INT7_STATUS_CORE0_CH3_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH3_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH3_INT7_STAT_BIT_OFFSET = 3;
  localparam int INT7_STATUS_CORE0_CH4_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH4_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH4_INT7_STAT_BIT_OFFSET = 4;
  localparam int INT7_STATUS_CORE0_CH5_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH5_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH5_INT7_STAT_BIT_OFFSET = 5;
  localparam int INT7_STATUS_CORE0_CH6_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH6_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH6_INT7_STAT_BIT_OFFSET = 6;
  localparam int INT7_STATUS_CORE0_CH7_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE0_CH7_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE0_CH7_INT7_STAT_BIT_OFFSET = 7;
  localparam int INT7_STATUS_CORE1_CH0_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH0_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH0_INT7_STAT_BIT_OFFSET = 8;
  localparam int INT7_STATUS_CORE1_CH1_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH1_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH1_INT7_STAT_BIT_OFFSET = 9;
  localparam int INT7_STATUS_CORE1_CH2_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH2_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH2_INT7_STAT_BIT_OFFSET = 10;
  localparam int INT7_STATUS_CORE1_CH3_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH3_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH3_INT7_STAT_BIT_OFFSET = 11;
  localparam int INT7_STATUS_CORE1_CH4_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH4_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH4_INT7_STAT_BIT_OFFSET = 12;
  localparam int INT7_STATUS_CORE1_CH5_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH5_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH5_INT7_STAT_BIT_OFFSET = 13;
  localparam int INT7_STATUS_CORE1_CH6_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH6_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH6_INT7_STAT_BIT_OFFSET = 14;
  localparam int INT7_STATUS_CORE1_CH7_INT7_STAT_BIT_WIDTH = 1;
  localparam bit INT7_STATUS_CORE1_CH7_INT7_STAT_BIT_MASK = 1'h1;
  localparam int INT7_STATUS_CORE1_CH7_INT7_STAT_BIT_OFFSET = 15;
  localparam int CORE0_JOINT_MODE_BYTE_WIDTH = 4;
  localparam int CORE0_JOINT_MODE_BYTE_SIZE = 4;
  localparam bit [12:0] CORE0_JOINT_MODE_BYTE_OFFSET = 13'h1030;
  localparam int CORE0_JOINT_MODE_CORE0_JOINT_MODE_BIT_WIDTH = 1;
  localparam bit CORE0_JOINT_MODE_CORE0_JOINT_MODE_BIT_MASK = 1'h1;
  localparam int CORE0_JOINT_MODE_CORE0_JOINT_MODE_BIT_OFFSET = 0;
  localparam int CORE1_JOINT_MODE_BYTE_WIDTH = 4;
  localparam int CORE1_JOINT_MODE_BYTE_SIZE = 4;
  localparam bit [12:0] CORE1_JOINT_MODE_BYTE_OFFSET = 13'h1034;
  localparam int CORE1_JOINT_MODE_CORE1_JOINT_MODE_BIT_WIDTH = 1;
  localparam bit CORE1_JOINT_MODE_CORE1_JOINT_MODE_BIT_MASK = 1'h1;
  localparam int CORE1_JOINT_MODE_CORE1_JOINT_MODE_BIT_OFFSET = 0;
  localparam int CORE0_PRIORITY_BYTE_WIDTH = 4;
  localparam int CORE0_PRIORITY_BYTE_SIZE = 4;
  localparam bit [12:0] CORE0_PRIORITY_BYTE_OFFSET = 13'h1038;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_TOP_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE0_PRIORITY_CORE0_RD_PRIO_TOP_NUM_BIT_MASK = 3'h7;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_TOP_NUM_BIT_OFFSET = 0;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_TOP_BIT_WIDTH = 1;
  localparam bit CORE0_PRIORITY_CORE0_RD_PRIO_TOP_BIT_MASK = 1'h1;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_TOP_BIT_OFFSET = 3;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_NUM_BIT_MASK = 3'h7;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_NUM_BIT_OFFSET = 4;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_BIT_WIDTH = 1;
  localparam bit CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_BIT_MASK = 1'h1;
  localparam int CORE0_PRIORITY_CORE0_RD_PRIO_HIGH_BIT_OFFSET = 7;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_TOP_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE0_PRIORITY_CORE0_WR_PRIO_TOP_NUM_BIT_MASK = 3'h7;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_TOP_NUM_BIT_OFFSET = 8;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_TOP_BIT_WIDTH = 1;
  localparam bit CORE0_PRIORITY_CORE0_WR_PRIO_TOP_BIT_MASK = 1'h1;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_TOP_BIT_OFFSET = 11;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_NUM_BIT_MASK = 3'h7;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_NUM_BIT_OFFSET = 12;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_BIT_WIDTH = 1;
  localparam bit CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_BIT_MASK = 1'h1;
  localparam int CORE0_PRIORITY_CORE0_WR_PRIO_HIGH_BIT_OFFSET = 15;
  localparam int CORE1_PRIORITY_BYTE_WIDTH = 4;
  localparam int CORE1_PRIORITY_BYTE_SIZE = 4;
  localparam bit [12:0] CORE1_PRIORITY_BYTE_OFFSET = 13'h103c;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_TOP_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE1_PRIORITY_CORE1_RD_PRIO_TOP_NUM_BIT_MASK = 3'h7;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_TOP_NUM_BIT_OFFSET = 0;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_TOP_BIT_WIDTH = 1;
  localparam bit CORE1_PRIORITY_CORE1_RD_PRIO_TOP_BIT_MASK = 1'h1;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_TOP_BIT_OFFSET = 3;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_NUM_BIT_MASK = 3'h7;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_NUM_BIT_OFFSET = 4;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_BIT_WIDTH = 1;
  localparam bit CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_BIT_MASK = 1'h1;
  localparam int CORE1_PRIORITY_CORE1_RD_PRIO_HIGH_BIT_OFFSET = 7;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_TOP_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE1_PRIORITY_CORE1_WR_PRIO_TOP_NUM_BIT_MASK = 3'h7;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_TOP_NUM_BIT_OFFSET = 8;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_TOP_BIT_WIDTH = 1;
  localparam bit CORE1_PRIORITY_CORE1_WR_PRIO_TOP_BIT_MASK = 1'h1;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_TOP_BIT_OFFSET = 11;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_NUM_BIT_WIDTH = 3;
  localparam bit [2:0] CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_NUM_BIT_MASK = 3'h7;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_NUM_BIT_OFFSET = 12;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_BIT_WIDTH = 1;
  localparam bit CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_BIT_MASK = 1'h1;
  localparam int CORE1_PRIORITY_CORE1_WR_PRIO_HIGH_BIT_OFFSET = 15;
  localparam int CORE0_CLKDIV_BYTE_WIDTH = 4;
  localparam int CORE0_CLKDIV_BYTE_SIZE = 4;
  localparam bit [12:0] CORE0_CLKDIV_BYTE_OFFSET = 13'h1040;
  localparam int CORE0_CLKDIV_CORE0_CLKDIV_RATIO_BIT_WIDTH = 4;
  localparam bit [3:0] CORE0_CLKDIV_CORE0_CLKDIV_RATIO_BIT_MASK = 4'hf;
  localparam int CORE0_CLKDIV_CORE0_CLKDIV_RATIO_BIT_OFFSET = 0;
  localparam int CORE1_CLKDIV_BYTE_WIDTH = 4;
  localparam int CORE1_CLKDIV_BYTE_SIZE = 4;
  localparam bit [12:0] CORE1_CLKDIV_BYTE_OFFSET = 13'h1044;
  localparam int CORE1_CLKDIV_CORE1_CLKDIV_RATIO_BIT_WIDTH = 4;
  localparam bit [3:0] CORE1_CLKDIV_CORE1_CLKDIV_RATIO_BIT_MASK = 4'hf;
  localparam int CORE1_CLKDIV_CORE1_CLKDIV_RATIO_BIT_OFFSET = 0;
  localparam int CORE0_CH_START_BYTE_WIDTH = 4;
  localparam int CORE0_CH_START_BYTE_SIZE = 4;
  localparam bit [12:0] CORE0_CH_START_BYTE_OFFSET = 13'h1048;
  localparam int CORE0_CH_START_CORE0_CHANNEL_START_BIT_WIDTH = 8;
  localparam bit [7:0] CORE0_CH_START_CORE0_CHANNEL_START_BIT_MASK = 8'hff;
  localparam int CORE0_CH_START_CORE0_CHANNEL_START_BIT_OFFSET = 0;
  localparam int CORE1_CH_START_BYTE_WIDTH = 4;
  localparam int CORE1_CH_START_BYTE_SIZE = 4;
  localparam bit [12:0] CORE1_CH_START_BYTE_OFFSET = 13'h104c;
  localparam int CORE1_CH_START_CORE1_CHANNEL_START_BIT_WIDTH = 8;
  localparam bit [7:0] CORE1_CH_START_CORE1_CHANNEL_START_BIT_MASK = 8'hff;
  localparam int CORE1_CH_START_CORE1_CHANNEL_START_BIT_OFFSET = 0;
  localparam int PERIPH_RX_CTRL_BYTE_WIDTH = 4;
  localparam int PERIPH_RX_CTRL_BYTE_SIZE = 4;
  localparam bit [12:0] PERIPH_RX_CTRL_BYTE_OFFSET = 13'h1050;
  localparam int PERIPH_RX_CTRL_PERIPH_RX_REQ_BIT_WIDTH = 31;
  localparam bit [30:0] PERIPH_RX_CTRL_PERIPH_RX_REQ_BIT_MASK = 31'h7fffffff;
  localparam int PERIPH_RX_CTRL_PERIPH_RX_REQ_BIT_OFFSET = 1;
  localparam int PERIPH_TX_CTRL_BYTE_WIDTH = 4;
  localparam int PERIPH_TX_CTRL_BYTE_SIZE = 4;
  localparam bit [12:0] PERIPH_TX_CTRL_BYTE_OFFSET = 13'h1054;
  localparam int PERIPH_TX_CTRL_PERIPH_TX_REQ_BIT_WIDTH = 31;
  localparam bit [30:0] PERIPH_TX_CTRL_PERIPH_TX_REQ_BIT_MASK = 31'h7fffffff;
  localparam int PERIPH_TX_CTRL_PERIPH_TX_REQ_BIT_OFFSET = 1;
  localparam int IDLE_BYTE_WIDTH = 4;
  localparam int IDLE_BYTE_SIZE = 4;
  localparam bit [12:0] IDLE_BYTE_OFFSET = 13'h10d0;
  localparam int IDLE_IDLE_BIT_WIDTH = 1;
  localparam bit IDLE_IDLE_BIT_MASK = 1'h1;
  localparam int IDLE_IDLE_BIT_OFFSET = 0;
  localparam int USER_DEF_STATUS_BYTE_WIDTH = 4;
  localparam int USER_DEF_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] USER_DEF_STATUS_BYTE_OFFSET = 13'h10e0;
  localparam int USER_DEF_STATUS_USER_DEF_INT_NUM_BIT_WIDTH = 4;
  localparam bit [3:0] USER_DEF_STATUS_USER_DEF_INT_NUM_BIT_MASK = 4'hf;
  localparam int USER_DEF_STATUS_USER_DEF_INT_NUM_BIT_OFFSET = 0;
  localparam int USER_DEF_STATUS_USER_DEF_DUAL_CORE_BIT_WIDTH = 1;
  localparam bit USER_DEF_STATUS_USER_DEF_DUAL_CORE_BIT_MASK = 1'h1;
  localparam int USER_DEF_STATUS_USER_DEF_DUAL_CORE_BIT_OFFSET = 5;
  localparam int USER_DEF_STATUS_USER_DEF_IC_BIT_WIDTH = 1;
  localparam bit USER_DEF_STATUS_USER_DEF_IC_BIT_MASK = 1'h1;
  localparam int USER_DEF_STATUS_USER_DEF_IC_BIT_OFFSET = 6;
  localparam int USER_DEF_STATUS_USER_DEF_IC_DUAL_PORT_BIT_WIDTH = 1;
  localparam bit USER_DEF_STATUS_USER_DEF_IC_DUAL_PORT_BIT_MASK = 1'h1;
  localparam int USER_DEF_STATUS_USER_DEF_IC_DUAL_PORT_BIT_OFFSET = 7;
  localparam int USER_DEF_STATUS_USER_DEF_CLKGATE_BIT_WIDTH = 1;
  localparam bit USER_DEF_STATUS_USER_DEF_CLKGATE_BIT_MASK = 1'h1;
  localparam int USER_DEF_STATUS_USER_DEF_CLKGATE_BIT_OFFSET = 8;
  localparam int USER_CORE0_DEF_STATUS0_BYTE_WIDTH = 4;
  localparam int USER_CORE0_DEF_STATUS0_BYTE_SIZE = 4;
  localparam bit [12:0] USER_CORE0_DEF_STATUS0_BYTE_OFFSET = 13'h10f0;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_CH_NUM_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_CH_NUM_BIT_MASK = 4'hf;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_CH_NUM_BIT_OFFSET = 0;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_FIFO_SIZE_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_FIFO_SIZE_BIT_MASK = 4'hf;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_FIFO_SIZE_BIT_OFFSET = 4;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_WCMD_DEPTH_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_WCMD_DEPTH_BIT_MASK = 4'hf;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_WCMD_DEPTH_BIT_OFFSET = 8;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_RCMD_DEPTH_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_RCMD_DEPTH_BIT_MASK = 4'hf;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_RCMD_DEPTH_BIT_OFFSET = 12;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_ADDR_BITS_BIT_WIDTH = 6;
  localparam bit [5:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_ADDR_BITS_BIT_MASK = 6'h3f;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_ADDR_BITS_BIT_OFFSET = 16;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_AXI_32_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_AXI_32_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_AXI_32_BIT_OFFSET = 22;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_BUFF_BITS_BIT_WIDTH = 5;
  localparam bit [4:0] USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_BUFF_BITS_BIT_MASK = 5'h1f;
  localparam int USER_CORE0_DEF_STATUS0_USER_DEF_CORE0_BUFF_BITS_BIT_OFFSET = 24;
  localparam int USER_CORE0_DEF_STATUS1_BYTE_WIDTH = 4;
  localparam int USER_CORE0_DEF_STATUS1_BYTE_SIZE = 4;
  localparam bit [12:0] USER_CORE0_DEF_STATUS1_BYTE_OFFSET = 13'h10f4;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WDT_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WDT_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WDT_BIT_OFFSET = 0;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TIMEOUT_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TIMEOUT_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TIMEOUT_BIT_OFFSET = 1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TOKENS_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TOKENS_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_TOKENS_BIT_OFFSET = 2;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PRIO_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PRIO_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PRIO_BIT_OFFSET = 3;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_OUTS_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_OUTS_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_OUTS_BIT_OFFSET = 4;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WAIT_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WAIT_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_WAIT_BIT_OFFSET = 5;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_BLOCK_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_BLOCK_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_BLOCK_BIT_OFFSET = 6;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_JOINT_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_JOINT_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_JOINT_BIT_OFFSET = 7;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_INDEPENDENT_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_INDEPENDENT_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_INDEPENDENT_BIT_OFFSET = 8;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PERIPH_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PERIPH_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_PERIPH_BIT_OFFSET = 9;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_LISTS_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_LISTS_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_LISTS_BIT_OFFSET = 10;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_END_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_END_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_END_BIT_OFFSET = 11;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_CLKDIV_BIT_WIDTH = 1;
  localparam bit USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_CLKDIV_BIT_MASK = 1'h1;
  localparam int USER_CORE0_DEF_STATUS1_USER_DEF_CORE0_CLKDIV_BIT_OFFSET = 12;
  localparam int USER_CORE1_DEF_STATUS0_BYTE_WIDTH = 4;
  localparam int USER_CORE1_DEF_STATUS0_BYTE_SIZE = 4;
  localparam bit [12:0] USER_CORE1_DEF_STATUS0_BYTE_OFFSET = 13'h10f8;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_CH_NUM_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_CH_NUM_BIT_MASK = 4'hf;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_CH_NUM_BIT_OFFSET = 0;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_FIFO_SIZE_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_FIFO_SIZE_BIT_MASK = 4'hf;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_FIFO_SIZE_BIT_OFFSET = 4;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_WCMD_DEPTH_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_WCMD_DEPTH_BIT_MASK = 4'hf;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_WCMD_DEPTH_BIT_OFFSET = 8;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_RCMD_DEPTH_BIT_WIDTH = 4;
  localparam bit [3:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_RCMD_DEPTH_BIT_MASK = 4'hf;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_RCMD_DEPTH_BIT_OFFSET = 12;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_ADDR_BITS_BIT_WIDTH = 6;
  localparam bit [5:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_ADDR_BITS_BIT_MASK = 6'h3f;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_ADDR_BITS_BIT_OFFSET = 16;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_AXI_32_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_AXI_32_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_AXI_32_BIT_OFFSET = 22;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_BUFF_BITS_BIT_WIDTH = 5;
  localparam bit [4:0] USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_BUFF_BITS_BIT_MASK = 5'h1f;
  localparam int USER_CORE1_DEF_STATUS0_USER_DEF_CORE1_BUFF_BITS_BIT_OFFSET = 24;
  localparam int USER_CORE1_DEF_STATUS1_BYTE_WIDTH = 4;
  localparam int USER_CORE1_DEF_STATUS1_BYTE_SIZE = 4;
  localparam bit [12:0] USER_CORE1_DEF_STATUS1_BYTE_OFFSET = 13'h10fc;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WDT_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WDT_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WDT_BIT_OFFSET = 0;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TIMEOUT_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TIMEOUT_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TIMEOUT_BIT_OFFSET = 1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TOKENS_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TOKENS_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_TOKENS_BIT_OFFSET = 2;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PRIO_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PRIO_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PRIO_BIT_OFFSET = 3;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_OUTS_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_OUTS_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_OUTS_BIT_OFFSET = 4;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WAIT_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WAIT_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_WAIT_BIT_OFFSET = 5;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_BLOCK_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_BLOCK_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_BLOCK_BIT_OFFSET = 6;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_JOINT_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_JOINT_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_JOINT_BIT_OFFSET = 7;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_INDEPENDENT_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_INDEPENDENT_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_INDEPENDENT_BIT_OFFSET = 8;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PERIPH_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PERIPH_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_PERIPH_BIT_OFFSET = 9;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_LISTS_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_LISTS_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_LISTS_BIT_OFFSET = 10;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_END_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_END_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_END_BIT_OFFSET = 11;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_CLKDIV_BIT_WIDTH = 1;
  localparam bit USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_CLKDIV_BIT_MASK = 1'h1;
  localparam int USER_CORE1_DEF_STATUS1_USER_DEF_CORE1_CLKDIV_BIT_OFFSET = 12;
endpackage
