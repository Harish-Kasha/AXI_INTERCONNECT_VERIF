`ifndef RAL_EXAMPLE_REG_BLOCK
`define RAL_EXAMPLE_REG_BLOCK

import uvm_pkg::*;

class ral_reg_example_reg_block_REG1 extends uvm_reg;
	rand uvm_reg_field reg1_field;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   reg1_field: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_REG1");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.reg1_field = uvm_reg_field::type_id::create("reg1_field",,get_full_name());
      this.reg1_field.configure(this, 32, 0, "RW", 0, 32'hABBADEAD, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_REG1)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_REG1


class ral_reg_example_reg_block_REG3 extends uvm_reg;
	rand uvm_reg_field reg3_field;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   reg3_field: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_REG3");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.reg3_field = uvm_reg_field::type_id::create("reg3_field",,get_full_name());
      this.reg3_field.configure(this, 32, 0, "RW", 0, 32'h000000, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_REG3)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_REG3


class ral_reg_example_reg_block_REG2 extends uvm_reg;
	rand uvm_reg_field reg2_field1;
	rand uvm_reg_field reg2_field2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   reg2_field1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	   reg2_field2: coverpoint {m_data[31:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "example_reg_block_REG2");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.reg2_field1 = uvm_reg_field::type_id::create("reg2_field1",,get_full_name());
      this.reg2_field1.configure(this, 16, 0, "RW", 0, 0, 1, 0, 1);
      this.reg2_field2 = uvm_reg_field::type_id::create("reg2_field2",,get_full_name());
      this.reg2_field2.configure(this, 16, 16, "RW", 0, 0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_REG2)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_REG2


class ral_reg_example_reg_block_A0 extends uvm_reg;
	rand uvm_reg_field a0_f;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   a0_f: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_A0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.a0_f = uvm_reg_field::type_id::create("a0_f",,get_full_name());
      this.a0_f.configure(this, 32, 0, "RW", 0, 0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_A0)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_A0


class ral_reg_example_reg_block_A1 extends uvm_reg;
	rand uvm_reg_field a1_f;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   a1_f: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_A1");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.a1_f = uvm_reg_field::type_id::create("a1_f",,get_full_name());
      this.a1_f.configure(this, 32, 0, "RW", 0, 0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_A1)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_A1


class ral_reg_example_reg_block_A2 extends uvm_reg;
	rand uvm_reg_field a2_f;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   a2_f: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_A2");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.a2_f = uvm_reg_field::type_id::create("a2_f",,get_full_name());
      this.a2_f.configure(this, 32, 0, "RW", 0, 0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_A2)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_A2


class ral_reg_example_reg_block_A3 extends uvm_reg;
	rand uvm_reg_field a3_f;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   a3_f: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "example_reg_block_A3");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.a3_f = uvm_reg_field::type_id::create("a3_f",,get_full_name());
      this.a3_f.configure(this, 32, 0, "RW", 0, 0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_example_reg_block_A3)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_example_reg_block_A3


class ral_block_example_reg_block extends uvm_reg_block;
	rand ral_reg_example_reg_block_REG1 REG1;
	rand ral_reg_example_reg_block_REG3 REG3;
	rand ral_reg_example_reg_block_REG2 REG2;
	rand ral_reg_example_reg_block_A0 A0;
	rand ral_reg_example_reg_block_A1 A1;
	rand ral_reg_example_reg_block_A2 A2;
	rand ral_reg_example_reg_block_A3 A3;
   local uvm_reg_data_t m_offset;
	rand uvm_reg_field REG1_reg1_field;
	rand uvm_reg_field reg1_field;
	rand uvm_reg_field REG3_reg3_field;
	rand uvm_reg_field reg3_field;
	rand uvm_reg_field REG2_reg2_field1;
	rand uvm_reg_field reg2_field1;
	rand uvm_reg_field REG2_reg2_field2;
	rand uvm_reg_field reg2_field2;
	rand uvm_reg_field A0_a0_f;
	rand uvm_reg_field a0_f;
	rand uvm_reg_field A1_a1_f;
	rand uvm_reg_field a1_f;
	rand uvm_reg_field A2_a2_f;
	rand uvm_reg_field a2_f;
	rand uvm_reg_field A3_a3_f;
	rand uvm_reg_field a3_f;


covergroup cg_addr (input string name);
	option.per_instance = 1;
option.name = get_name();

	REG1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h80000000 };
		option.weight = 1;
	}

	REG3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hACDCACDC };
		option.weight = 1;
	}

	REG2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h80000008 };
		option.weight = 1;
	}

	A0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h800 };
		option.weight = 1;
	}

	A1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h804 };
		option.weight = 1;
	}

	A2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h808 };
		option.weight = 1;
	}

	A3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h80C };
		option.weight = 1;
	}
endgroup
	function new(string name = "example_reg_block");
		super.new(name, build_coverage(UVM_CVR_ADDR_MAP));
		if (has_coverage(UVM_CVR_ADDR_MAP))
			cg_addr = new("cg_addr");
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 4, UVM_LITTLE_ENDIAN, 0);
      this.REG1 = ral_reg_example_reg_block_REG1::type_id::create("REG1",,get_full_name());
      if(this.REG1.has_coverage(UVM_CVR_REG_BITS))
      	this.REG1.cg_bits.option.name = "REG1";
      this.REG1.configure(this, null, "");
      this.REG1.build();
      this.default_map.add_reg(this.REG1, `UVM_REG_ADDR_WIDTH'h80000000, "RW", 0);
		this.REG1_reg1_field = this.REG1.reg1_field;
		this.reg1_field = this.REG1.reg1_field;
      this.REG3 = ral_reg_example_reg_block_REG3::type_id::create("REG3",,get_full_name());
      if(this.REG3.has_coverage(UVM_CVR_REG_BITS))
      	this.REG3.cg_bits.option.name = "REG3";
      this.REG3.configure(this, null, "");
      this.REG3.build();
      this.default_map.add_reg(this.REG3, `UVM_REG_ADDR_WIDTH'hACDCACDC, "RW", 0);
		this.REG3_reg3_field = this.REG3.reg3_field;
		this.reg3_field = this.REG3.reg3_field;
      this.REG2 = ral_reg_example_reg_block_REG2::type_id::create("REG2",,get_full_name());
      if(this.REG2.has_coverage(UVM_CVR_REG_BITS))
      	this.REG2.cg_bits.option.name = "REG2";
      this.REG2.configure(this, null, "");
      this.REG2.build();
      this.default_map.add_reg(this.REG2, `UVM_REG_ADDR_WIDTH'h80000008, "RW", 0);
		this.REG2_reg2_field1 = this.REG2.reg2_field1;
		this.reg2_field1 = this.REG2.reg2_field1;
		this.REG2_reg2_field2 = this.REG2.reg2_field2;
		this.reg2_field2 = this.REG2.reg2_field2;
      this.A0 = ral_reg_example_reg_block_A0::type_id::create("A0",,get_full_name());
      if(this.A0.has_coverage(UVM_CVR_REG_BITS))
      	this.A0.cg_bits.option.name = "A0";
      this.A0.configure(this, null, "");
      this.A0.build();
      this.default_map.add_reg(this.A0, `UVM_REG_ADDR_WIDTH'h800, "RW", 0);
		this.A0_a0_f = this.A0.a0_f;
		this.a0_f = this.A0.a0_f;
      this.A1 = ral_reg_example_reg_block_A1::type_id::create("A1",,get_full_name());
      if(this.A1.has_coverage(UVM_CVR_REG_BITS))
      	this.A1.cg_bits.option.name = "A1";
      this.A1.configure(this, null, "");
      this.A1.build();
      this.default_map.add_reg(this.A1, `UVM_REG_ADDR_WIDTH'h804, "RW", 0);
		this.A1_a1_f = this.A1.a1_f;
		this.a1_f = this.A1.a1_f;
      this.A2 = ral_reg_example_reg_block_A2::type_id::create("A2",,get_full_name());
      if(this.A2.has_coverage(UVM_CVR_REG_BITS))
      	this.A2.cg_bits.option.name = "A2";
      this.A2.configure(this, null, "");
      this.A2.build();
      this.default_map.add_reg(this.A2, `UVM_REG_ADDR_WIDTH'h808, "RW", 0);
		this.A2_a2_f = this.A2.a2_f;
		this.a2_f = this.A2.a2_f;
      this.A3 = ral_reg_example_reg_block_A3::type_id::create("A3",,get_full_name());
      if(this.A3.has_coverage(UVM_CVR_REG_BITS))
      	this.A3.cg_bits.option.name = "A3";
      this.A3.configure(this, null, "");
      this.A3.build();
      this.default_map.add_reg(this.A3, `UVM_REG_ADDR_WIDTH'h80C, "RW", 0);
		this.A3_a3_f = this.A3.a3_f;
		this.a3_f = this.A3.a3_f;
   endfunction : build

	`uvm_object_utils(ral_block_example_reg_block)


function void sample(uvm_reg_addr_t offset,
                     bit            is_read,
                     uvm_reg_map    map);
  if (get_coverage(UVM_CVR_ADDR_MAP)) begin
    m_offset = offset;
    cg_addr.sample();
  end
endfunction
endclass : ral_block_example_reg_block



`endif

